module dff_from_nand();
wire Q,Q_BAR;
reg D,CLK;
nand U1 (X,D,CLK) ;
nand U2 (Y,X,CLK) ;
nand U3 (Q,Q_BAR,X);
nand U4 (Q_BAR,Q,Y);
// Testbench of above code
 initial begin
 $monitor ( "CLK = %b D = %b Q = %b Q_BAR = %b" ,CLK, D, Q, Q_BAR);
 CLK = 0;
 D = 0;
 #3 D = 1;
 #3 D = 0;
 #3 $finish ;
 end
 always #2 CLK = ~CLK;

 endmodule